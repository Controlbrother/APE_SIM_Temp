<?xml version="1.0" encoding="UTF-8" standalone="no"?>
<Root>
	<creator type="key">ConfigurationDesk 6.6</creator>
	<application>
		<Name type="key">NoaApp.CDL</Name>
		<DisplayName type="key">NoaApp</DisplayName>
		<Path type="key">.\NoaApp</Path>
		<Component type="key">ProjectApplication</Component>
		<Type type="key">14</Type>
		<ApplicationType type="key">3</ApplicationType>
		<Flags type="key">41216</Flags>
		<ItemInfoDate type="key">2021/6/8 11:23:30</ItemInfoDate>
		<ItemInfoPath type="key">$FPATH$</ItemInfoPath>
		<ItemInfoDocs type="key"/>
		<ItemInfoDescr type="key"/>
		<ItemInfoAuthor type="key">Cheng</ItemInfoAuthor>
		<Log type="key"/>
		<AddInfoDb type="key"/>
		<DatabaseID type="key">-1</DatabaseID>
		<EntityID type="key">{25B58803-3EFF-4AAD-96D5-DEF59FA3602A}</EntityID>
		<item>
			<Name type="key">WindowConfiguration.xml</Name>
			<DisplayName type="key">WindowConfiguration.xml</DisplayName>
			<Path type="key">.</Path>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">260</Flags>
			<ExtendedFlags type="key">16</ExtendedFlags>
			<Type type="key">4</Type>
			<ItemInfoDate type="key">2020/8/8 10:58:43</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">GW00216231</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{8A2B69BE-B703-44D9-A9AD-33B753E4F195}</EntityID>
			<Targets/>
		</item>
		<item>
			<DisplayName type="key">Device Topology</DisplayName>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">131328</Flags>
			<ExtendedFlags type="key">16</ExtendedFlags>
			<Type type="key">33</Type>
			<ItemInfoDate type="key">2020/8/8 10:58:43</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">GW00216231</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{F898C2BC-52A9-4748-BFB4-963D5D2268C7}</EntityID>
			<Targets/>
		</item>
		<item>
			<DisplayName type="key">Hardware Topology</DisplayName>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">256</Flags>
			<ExtendedFlags type="key">16</ExtendedFlags>
			<Type type="key">19</Type>
			<ItemInfoDate type="key">2020/8/8 10:58:43</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">GW00216231</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{45CF0532-6B5F-4DEB-A0BA-122548B320B4}</EntityID>
			<Targets/>
		</item>
		<item>
			<DisplayName type="key">Model Topology</DisplayName>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">256</Flags>
			<ExtendedFlags type="key">16</ExtendedFlags>
			<Type type="key">31</Type>
			<ItemInfoDate type="key">2020/8/8 10:58:43</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">GW00216231</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key">Model location:
F:\05_dspace_Work_Files\11_HWA_Project\Git_ADAS_Store\projcct\adas_project\Noa_Nofusion.slx
</Log>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{FABCC1B7-F34C-4A0E-8657-FF02FD24149A}</EntityID>
			<Targets/>
		</item>
		<item>
			<DisplayName type="key">Communication Matrices</DisplayName>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">256</Flags>
			<ExtendedFlags type="key">16</ExtendedFlags>
			<Type type="key">70</Type>
			<ItemInfoDate type="key">2020/8/8 10:58:43</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">GW00216231</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{02903D02-F798-4922-B7E4-A804BBE0EDF7}</EntityID>
			<Targets/>
		</item>
		<item>
			<DisplayName type="key">External Cable Harness</DisplayName>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">131328</Flags>
			<ExtendedFlags type="key">16</ExtendedFlags>
			<Type type="key">32</Type>
			<ItemInfoDate type="key">2020/8/8 10:58:43</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">GW00216231</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{BDD70D61-CB95-438E-BC39-D669A73035F4}</EntityID>
			<Targets/>
		</item>
		<item>
			<Name type="key">Application.cfgx</Name>
			<DisplayName type="key">Core Application</DisplayName>
			<Path type="key">.</Path>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">260</Flags>
			<ExtendedFlags type="key">16</ExtendedFlags>
			<Type type="key">20</Type>
			<ItemInfoDate type="key">2020/8/8 10:58:43</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">GW00216231</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{768A4438-04CF-4B37-98A7-043AF737ADBF}</EntityID>
			<Targets/>
		</item>
		<item>
			<Name type="key">Build Results</Name>
			<DisplayName type="key">Build Results</DisplayName>
			<Path type="key">.</Path>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">256</Flags>
			<ExtendedFlags type="key">0</ExtendedFlags>
			<Type type="key">58</Type>
			<ItemInfoDate type="key">2021/8/4 10:29:35</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">GW00216231</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{C7DF596A-E104-406F-BFC5-0E4FF02BF0C2}</EntityID>
			<Targets/>
			<item>
				<Name type="key">Build Results</Name>
				<DisplayName type="key">Noa_Nofusion</DisplayName>
				<Path type="key">.</Path>
				<Component type="key">ProjectApplication</Component>
				<Flags type="key">260</Flags>
				<ExtendedFlags type="key">0</ExtendedFlags>
				<Type type="key">29</Type>
				<ItemInfoDate type="key">2021/8/31 11:13:43</ItemInfoDate>
				<ItemInfoPath type="key"/>
				<ItemInfoDocs type="key"/>
				<ItemInfoDescr type="key"/>
				<ItemInfoAuthor type="key">GW00216231</ItemInfoAuthor>
				<ItemInfoAddInfoDb type="key"/>
				<Log type="key"/>
				<DatabaseID type="key">-1</DatabaseID>
				<EntityID type="key">{EBBB3943-7F6F-463D-8ADF-78DBE0D5F8CA}</EntityID>
				<Targets/>
				<item>
					<Name type="key">Noa_Nofusion.a2l</Name>
					<DisplayName type="key">Noa_Nofusion.a2l</DisplayName>
					<Path type="key">.\Build Results</Path>
					<Component type="key">ProjectApplication</Component>
					<Flags type="key">256</Flags>
					<ExtendedFlags type="key">0</ExtendedFlags>
					<Type type="key">60</Type>
					<ItemInfoDate type="key">2021/8/31 11:13:43</ItemInfoDate>
					<ItemInfoPath type="key"/>
					<ItemInfoDocs type="key"/>
					<ItemInfoDescr type="key"/>
					<ItemInfoAuthor type="key">GW00216231</ItemInfoAuthor>
					<ItemInfoAddInfoDb type="key"/>
					<Log type="key"/>
					<DatabaseID type="key">-1</DatabaseID>
					<EntityID type="key">{E9FA17F7-97C4-48F4-B8D8-01015EED3A2A}</EntityID>
					<Targets/>
				</item>
			</item>
			<item>
				<Name type="key">Build Results</Name>
				<DisplayName type="key">itSDFROOT</DisplayName>
				<Path type="key">.</Path>
				<Component type="key">ProjectApplication</Component>
				<Flags type="key">260</Flags>
				<ExtendedFlags type="key">0</ExtendedFlags>
				<Type type="key">29</Type>
				<ItemInfoDate type="key">2021/8/4 10:29:35</ItemInfoDate>
				<ItemInfoPath type="key"/>
				<ItemInfoDocs type="key"/>
				<ItemInfoDescr type="key"/>
				<ItemInfoAuthor type="key">GW00216231</ItemInfoAuthor>
				<ItemInfoAddInfoDb type="key"/>
				<Log type="key"/>
				<DatabaseID type="key">-1</DatabaseID>
				<EntityID type="key">{B1777828-A282-42B0-9DBE-589DC718C3C4}</EntityID>
				<Targets/>
				<item>
					<Name type="key">Noa_Nofusion.expswcfg</Name>
					<DisplayName type="key">Noa_Nofusion.expswcfg</DisplayName>
					<Path type="key">.\Build Results</Path>
					<Component type="key">ProjectApplication</Component>
					<Flags type="key">256</Flags>
					<ExtendedFlags type="key">0</ExtendedFlags>
					<Type type="key">71</Type>
					<ItemInfoDate type="key">2021/8/4 10:29:35</ItemInfoDate>
					<ItemInfoPath type="key"/>
					<ItemInfoDocs type="key"/>
					<ItemInfoDescr type="key"/>
					<ItemInfoAuthor type="key">GW00216231</ItemInfoAuthor>
					<ItemInfoAddInfoDb type="key"/>
					<Log type="key"/>
					<DatabaseID type="key">-1</DatabaseID>
					<EntityID type="key">{F972570E-C47C-46AB-9D3E-54EF79E05BB4}</EntityID>
					<Targets/>
				</item>
				<item>
					<Name type="key">Noa_Nofusion.map</Name>
					<DisplayName type="key">Noa_Nofusion.map</DisplayName>
					<Path type="key">.\Build Results</Path>
					<Component type="key">ProjectApplication</Component>
					<Flags type="key">256</Flags>
					<ExtendedFlags type="key">0</ExtendedFlags>
					<Type type="key">36</Type>
					<ItemInfoDate type="key">2021/8/4 10:29:35</ItemInfoDate>
					<ItemInfoPath type="key"/>
					<ItemInfoDocs type="key"/>
					<ItemInfoDescr type="key"/>
					<ItemInfoAuthor type="key">GW00216231</ItemInfoAuthor>
					<ItemInfoAddInfoDb type="key"/>
					<Log type="key"/>
					<DatabaseID type="key">-1</DatabaseID>
					<EntityID type="key">{6900B0D9-CEEF-4528-95DA-1349D39828F4}</EntityID>
					<Targets/>
				</item>
				<item>
					<Name type="key">Noa_Nofusion.s19</Name>
					<DisplayName type="key">Noa_Nofusion.s19</DisplayName>
					<Path type="key">.\Build Results</Path>
					<Component type="key">ProjectApplication</Component>
					<Flags type="key">256</Flags>
					<ExtendedFlags type="key">0</ExtendedFlags>
					<Type type="key">36</Type>
					<ItemInfoDate type="key">2021/8/31 11:13:43</ItemInfoDate>
					<ItemInfoPath type="key"/>
					<ItemInfoDocs type="key"/>
					<ItemInfoDescr type="key"/>
					<ItemInfoAuthor type="key">GW00216231</ItemInfoAuthor>
					<ItemInfoAddInfoDb type="key"/>
					<Log type="key"/>
					<DatabaseID type="key">-1</DatabaseID>
					<EntityID type="key">{0A161E8D-5C3D-4286-B5FE-CF146871F1B7}</EntityID>
					<Targets/>
				</item>
				<item>
					<Name type="key">Noa_Nofusion.trc</Name>
					<DisplayName type="key">Noa_Nofusion.trc</DisplayName>
					<Path type="key">.\Build Results</Path>
					<Component type="key">ProjectApplication</Component>
					<Flags type="key">256</Flags>
					<ExtendedFlags type="key">0</ExtendedFlags>
					<Type type="key">34</Type>
					<ItemInfoDate type="key">2021/8/4 10:29:35</ItemInfoDate>
					<ItemInfoPath type="key"/>
					<ItemInfoDocs type="key"/>
					<ItemInfoDescr type="key"/>
					<ItemInfoAuthor type="key">GW00216231</ItemInfoAuthor>
					<ItemInfoAddInfoDb type="key"/>
					<Log type="key"/>
					<DatabaseID type="key">-1</DatabaseID>
					<EntityID type="key">{4EF01804-3344-4E43-A9FD-520353B075D3}</EntityID>
					<Targets/>
				</item>
				<item>
					<Name type="key">NoaApp.dsbuildinfo</Name>
					<DisplayName type="key">NoaApp.dsbuildinfo</DisplayName>
					<Path type="key">.\Build Results</Path>
					<Component type="key">ProjectApplication</Component>
					<Flags type="key">260</Flags>
					<ExtendedFlags type="key">0</ExtendedFlags>
					<Type type="key">4</Type>
					<ItemInfoDate type="key">2021/8/4 10:29:35</ItemInfoDate>
					<ItemInfoPath type="key"/>
					<ItemInfoDocs type="key"/>
					<ItemInfoDescr type="key"/>
					<ItemInfoAuthor type="key">GW00216231</ItemInfoAuthor>
					<ItemInfoAddInfoDb type="key"/>
					<Log type="key"/>
					<DatabaseID type="key">-1</DatabaseID>
					<EntityID type="key">{C83B9AAE-64F8-4613-8EC4-072C5F4CFBD6}</EntityID>
					<Targets/>
				</item>
				<item>
					<Name type="key">NoaApp.rta</Name>
					<DisplayName type="key">NoaApp.rta</DisplayName>
					<Path type="key">.\Build Results</Path>
					<Component type="key">ProjectApplication</Component>
					<Flags type="key">256</Flags>
					<ExtendedFlags type="key">0</ExtendedFlags>
					<Type type="key">37</Type>
					<ItemInfoDate type="key">2021/8/4 10:29:35</ItemInfoDate>
					<ItemInfoPath type="key"/>
					<ItemInfoDocs type="key"/>
					<ItemInfoDescr type="key"/>
					<ItemInfoAuthor type="key">GW00216231</ItemInfoAuthor>
					<ItemInfoAddInfoDb type="key"/>
					<Log type="key"/>
					<DatabaseID type="key">-1</DatabaseID>
					<EntityID type="key">{D1B6CF43-0CA6-475C-8952-D4E57419BBD6}</EntityID>
					<Targets/>
				</item>
				<item>
					<Name type="key">NoaApp.sdf</Name>
					<DisplayName type="key">NoaApp.sdf</DisplayName>
					<Path type="key">.\Build Results</Path>
					<Component type="key">ProjectApplication</Component>
					<Flags type="key">256</Flags>
					<ExtendedFlags type="key">0</ExtendedFlags>
					<Type type="key">35</Type>
					<ItemInfoDate type="key">2021/8/4 10:29:35</ItemInfoDate>
					<ItemInfoPath type="key"/>
					<ItemInfoDocs type="key"/>
					<ItemInfoDescr type="key"/>
					<ItemInfoAuthor type="key">GW00216231</ItemInfoAuthor>
					<ItemInfoAddInfoDb type="key"/>
					<Log type="key"/>
					<DatabaseID type="key">-1</DatabaseID>
					<EntityID type="key">{796B0A37-4D5F-4B48-9281-49C217367107}</EntityID>
					<Targets/>
				</item>
			</item>
		</item>
	</application>
</Root>